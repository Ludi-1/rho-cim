-- VHDL package for custom datatype (2d vector)
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package cnn_package is
        type data_array is array(natural range <>) of std_logic_vector;
end package;