module mlp_l_d8_c128_top #(
	datatype_size = 8,
	xbar_size = 128,
	output_datatype_size = 8
) (
input clk,
input rst
);
endmodule