module cnn_2_d2_c256_top #(
	datatype_size = 2,
	xbar_size = 256,
	output_datatype_size = 2
) (
input clk,
input rst
);
endmodule