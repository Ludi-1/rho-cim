module mlp_l_d4_c256_top #(
	datatype_size = 4,
	xbar_size = 256,
	output_datatype_size = 4
) (
input clk,
input rst
);
endmodule