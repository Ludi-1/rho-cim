module mlp_m_d2_c128_top #(
	datatype_size = 2,
	xbar_size = 128,
	output_datatype_size = 2
) (
input clk,
input rst
);
endmodule