module mlp_m_d4_c128_top #(
	datatype_size = 4,
	xbar_size = 128,
	output_datatype_size = 4
) (
input clk,
input rst
);
endmodule