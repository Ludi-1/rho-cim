module cnn_1_d4_c512_top #(
	datatype_size = 4,
	xbar_size = 512,
	output_datatype_size = 4
) (
input clk,
input rst
);
endmodule