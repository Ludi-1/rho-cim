module mlp_s_d8_c256_top #(
	datatype_size = 8,
	xbar_size = 256,
	output_datatype_size = 8
) (
input clk,
input rst
);
endmodule