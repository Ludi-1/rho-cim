typedef enum {
  S0, // Reset
  S1, // Idle
  S2, // Busy
  S3 // Start next
} state;

module fc_ctrl #(
    parameter datatype_size = 8,
    parameter input_size = 201,
    parameter xbar_size = 256,
    parameter v_cim_tiles = (input_size + xbar_size - 1) / xbar_size // ceiled division
) (
    input clk,
    input rst,
    input i_start,
    input i_cim_busy,
    output reg o_cim_we,
    input i_func_busy,
    output reg o_busy,
    input [datatype_size-1:0] i_data,
    output reg [$clog2(input_size)-1:0] o_ibuf_addr,
    output reg [$clog2(xbar_size)-1:0] o_cim_addr,
    output reg [datatype_size-1:0] o_data [v_cim_tiles-1:0]
);

int unsigned cim_addr, next_cim_addr;
int unsigned input_count, next_input_count;
state ctrl_state, next_ctrl_state;

assign o_cim_addr = cim_addr[$clog2(xbar_size)-1:0];
assign o_ibuf_addr = input_count[$clog2(input_size)-1:0];

genvar i;
generate
    for (i = 0; i < v_cim_tiles; i++) begin
        assign o_data[i] = i_data;
    end
endgenerate

always_ff @(posedge clk) begin
    if (rst) begin
        ctrl_state = S0;
        input_count = 0;
        cim_addr = 0;
    end else begin
        ctrl_state = next_ctrl_state;
        input_count = next_input_count;
        cim_addr = next_cim_addr;
    end
end

always_comb begin
    case (ctrl_state)
        S0: begin // Reset state
            next_input_count = 0;
            next_cim_addr = 0;
            if (i_start & !rst) begin // Start signal comes in
                o_busy = 1;
                if (i_cim_busy) begin // If next module busy
                    next_ctrl_state = S1; // Idle until not busy
                end else begin // If next module not busy
                    next_ctrl_state = S2; // Start transfer
                end
            end else begin // Stay in reset state
                o_cim_we = 0;
                o_busy = 0;
                next_ctrl_state = S0;
            end
        end
        S1: begin // Idle state
            o_busy = 1;
            next_input_count = 0;
            next_cim_addr = 0;
            if (!i_cim_busy) begin
                o_cim_we = 1;
                next_ctrl_state = S2;
            end else begin
                o_cim_we = 0;
                next_ctrl_state = S1;
            end
        end
        S2: begin // Busy state
            o_busy = 1;
            if (input_count >= input_size - 1) begin
                o_cim_we = 0;
                if (!i_func_busy) begin
                    next_ctrl_state = S3; // Start
                    next_input_count = 0;
                    next_cim_addr = 0;
                end else begin
                    next_ctrl_state = S2;
                    next_input_count = input_count;
                    next_cim_addr = cim_addr;
                end
            end else begin
                o_cim_we = 1;
                next_ctrl_state = S2;
                next_input_count = input_count + 1;
                if (cim_addr >= xbar_size - 1) begin
                    next_cim_addr = 0;
                end else begin
                    next_cim_addr = cim_addr + 1;
                end
            end
        end
        S3: begin
            o_busy = 0;
            o_cim_we = 0;
            next_cim_addr = 0;
            next_input_count = 0;
            if (i_cim_busy) begin
                next_ctrl_state = S0;
            end else begin
                next_ctrl_state = S3;
            end
        end
        default: next_ctrl_state = S0;
    endcase
end

// `ifdef COCOTB_SIM
// initial begin
//     $dumpfile ("output/ibuf.fst");
//     for(int fifo_idx = 0; fifo_idx < fifo_length; fifo_idx ++) begin
//         $dumpvars (0, o_data[fifo_idx]);
//     end
//   #1;
// end
// `endif

endmodule
